module detector

// FIXME
const known_linkers = [
	// GNU ld
	// llvm-ld
	// link.exe
]