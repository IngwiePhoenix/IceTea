module detector

// FIXME
const known_archivers = [
	// GNU ar
	// llvm-ar
	// lib.exe
]