module detector

// FIXME
const known_archivers = []